module top_module(
    input clk,
    input areset,
    input j,
    input k,
    output out); 

    parameter OFF=1'b0, ON=1'b1; 
    reg state, next_state;

    always @(*) begin
        case (state)
            OFF:next_state=j?ON:OFF;
            ON:next_state=k?OFF:ON;
        endcase
    end
    always @(posedge clk, posedge areset) begin
        if(areset) state<=OFF;
        else state<=next_state;
    end
    assign out=(state==ON)?1'b1:1'b0;
endmodule
